
module clk_buf (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
